module CPU_top(
    
    );
endmodule